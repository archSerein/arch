module seg (data, seg1, seg0);
  
  input [7:0] data;
  output [6:0] seg1;
  output [6:0] seg0;

  assign seg0 = (data[3:0] == 4'b0000) ? 7'b0000001 :
                (data[3:0] == 4'b0001) ? 7'b1001111 :
                (data[3:0] == 4'b0010) ? 7'b0010010 :
                (data[3:0] == 4'b0011) ? 7'b0000110 :
                (data[3:0] == 4'b0100) ? 7'b1001100 :
                (data[3:0] == 4'b0101) ? 7'b0100100 :
                (data[3:0] == 4'b0110) ? 7'b0100000 :
                (data[3:0] == 4'b0111) ? 7'b0001111 :
                (data[3:0] == 4'b1000) ? 7'b0000000 :
                (data[3:0] == 4'b1001) ? 7'b0000100 :
                (data[3:0] == 4'b1010) ? 7'b0001000 :
                (data[3:0] == 4'b1011) ? 7'b1100000 :
                (data[3:0] == 4'b1100) ? 7'b0110001 :
                (data[3:0] == 4'b1101) ? 7'b1000010 :
                (data[3:0] == 4'b1110) ? 7'b0110000 :
                (data[3:0] == 4'b1111) ? 7'b0111000 :
                7'b1111111;


  assign seg1 = (data[7:4] == 4'b0000) ? 7'b0000001 :
                (data[7:4] == 4'b0001) ? 7'b1001111 :
                (data[7:4] == 4'b0010) ? 7'b0010010 :
                (data[7:4] == 4'b0011) ? 7'b0000110 :
                (data[7:4] == 4'b0100) ? 7'b1001100 :
                (data[7:4] == 4'b0101) ? 7'b0100100 :
                (data[7:4] == 4'b0110) ? 7'b0100000 :
                (data[7:4] == 4'b0111) ? 7'b0001111 :
                (data[7:4] == 4'b1000) ? 7'b0000000 :
                (data[7:4] == 4'b1001) ? 7'b0000100 :
                (data[7:4] == 4'b1010) ? 7'b0001000 :
                (data[7:4] == 4'b1011) ? 7'b1100000 :
                (data[7:4] == 4'b1100) ? 7'b0110001 :
                (data[7:4] == 4'b1101) ? 7'b1000010 :
                (data[7:4] == 4'b1110) ? 7'b0110000 :
                (data[7:4] == 4'b1111) ? 7'b0111000 :
                7'b1111111;

endmodule

