
module uart (
  output tx,
  input rx
);
  assign tx = rx;
endmodule
